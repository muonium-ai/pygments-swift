-- VHDL sample
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fib is
end entity;

architecture rtl of fib is
begin
  -- demo only
end architecture;
